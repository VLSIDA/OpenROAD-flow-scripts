VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram130_64x62
  FOREIGN fakeram130_64x62 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 189.980 BY 233.920 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 5.850 0.800 6.150 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 6.450 0.800 6.750 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 7.050 0.800 7.350 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 7.650 0.800 7.950 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 8.250 0.800 8.550 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 8.850 0.800 9.150 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 9.450 0.800 9.750 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 10.050 0.800 10.350 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 10.650 0.800 10.950 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 11.250 0.800 11.550 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 11.850 0.800 12.150 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 12.450 0.800 12.750 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 13.050 0.800 13.350 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 13.650 0.800 13.950 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 14.250 0.800 14.550 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 14.850 0.800 15.150 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 15.450 0.800 15.750 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 16.050 0.800 16.350 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 16.650 0.800 16.950 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 17.250 0.800 17.550 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 17.850 0.800 18.150 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 18.450 0.800 18.750 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 19.050 0.800 19.350 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 19.650 0.800 19.950 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 20.250 0.800 20.550 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 20.850 0.800 21.150 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 21.450 0.800 21.750 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 22.050 0.800 22.350 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 22.650 0.800 22.950 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 23.250 0.800 23.550 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 23.850 0.800 24.150 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 24.450 0.800 24.750 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 25.050 0.800 25.350 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 25.650 0.800 25.950 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 26.250 0.800 26.550 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 26.850 0.800 27.150 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 27.450 0.800 27.750 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 28.050 0.800 28.350 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 28.650 0.800 28.950 ;
    END
  END w_mask_in[38]
  PIN w_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 29.250 0.800 29.550 ;
    END
  END w_mask_in[39]
  PIN w_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 29.850 0.800 30.150 ;
    END
  END w_mask_in[40]
  PIN w_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 30.450 0.800 30.750 ;
    END
  END w_mask_in[41]
  PIN w_mask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 31.050 0.800 31.350 ;
    END
  END w_mask_in[42]
  PIN w_mask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 31.650 0.800 31.950 ;
    END
  END w_mask_in[43]
  PIN w_mask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 32.250 0.800 32.550 ;
    END
  END w_mask_in[44]
  PIN w_mask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 32.850 0.800 33.150 ;
    END
  END w_mask_in[45]
  PIN w_mask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 33.450 0.800 33.750 ;
    END
  END w_mask_in[46]
  PIN w_mask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 34.050 0.800 34.350 ;
    END
  END w_mask_in[47]
  PIN w_mask_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 34.650 0.800 34.950 ;
    END
  END w_mask_in[48]
  PIN w_mask_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 35.250 0.800 35.550 ;
    END
  END w_mask_in[49]
  PIN w_mask_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 35.850 0.800 36.150 ;
    END
  END w_mask_in[50]
  PIN w_mask_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 36.450 0.800 36.750 ;
    END
  END w_mask_in[51]
  PIN w_mask_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 37.050 0.800 37.350 ;
    END
  END w_mask_in[52]
  PIN w_mask_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 37.650 0.800 37.950 ;
    END
  END w_mask_in[53]
  PIN w_mask_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 38.250 0.800 38.550 ;
    END
  END w_mask_in[54]
  PIN w_mask_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 38.850 0.800 39.150 ;
    END
  END w_mask_in[55]
  PIN w_mask_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 39.450 0.800 39.750 ;
    END
  END w_mask_in[56]
  PIN w_mask_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 40.050 0.800 40.350 ;
    END
  END w_mask_in[57]
  PIN w_mask_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 40.650 0.800 40.950 ;
    END
  END w_mask_in[58]
  PIN w_mask_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 41.250 0.800 41.550 ;
    END
  END w_mask_in[59]
  PIN w_mask_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 41.850 0.800 42.150 ;
    END
  END w_mask_in[60]
  PIN w_mask_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 42.450 0.800 42.750 ;
    END
  END w_mask_in[61]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 68.250 0.800 68.550 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 68.850 0.800 69.150 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 69.450 0.800 69.750 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 70.050 0.800 70.350 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 70.650 0.800 70.950 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 71.250 0.800 71.550 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 71.850 0.800 72.150 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 72.450 0.800 72.750 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 73.050 0.800 73.350 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 73.650 0.800 73.950 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 74.250 0.800 74.550 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 74.850 0.800 75.150 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 75.450 0.800 75.750 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 76.050 0.800 76.350 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 76.650 0.800 76.950 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 77.250 0.800 77.550 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 77.850 0.800 78.150 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 78.450 0.800 78.750 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 79.050 0.800 79.350 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 79.650 0.800 79.950 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 80.250 0.800 80.550 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 80.850 0.800 81.150 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 81.450 0.800 81.750 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 82.050 0.800 82.350 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 82.650 0.800 82.950 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 83.250 0.800 83.550 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 83.850 0.800 84.150 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 84.450 0.800 84.750 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 85.050 0.800 85.350 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 85.650 0.800 85.950 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 86.250 0.800 86.550 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 86.850 0.800 87.150 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 87.450 0.800 87.750 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 88.050 0.800 88.350 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 88.650 0.800 88.950 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 89.250 0.800 89.550 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 89.850 0.800 90.150 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 90.450 0.800 90.750 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 91.050 0.800 91.350 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 91.650 0.800 91.950 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 92.250 0.800 92.550 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 92.850 0.800 93.150 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 93.450 0.800 93.750 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 94.050 0.800 94.350 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 94.650 0.800 94.950 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 95.250 0.800 95.550 ;
    END
  END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 95.850 0.800 96.150 ;
    END
  END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 96.450 0.800 96.750 ;
    END
  END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 97.050 0.800 97.350 ;
    END
  END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 97.650 0.800 97.950 ;
    END
  END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 98.250 0.800 98.550 ;
    END
  END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 98.850 0.800 99.150 ;
    END
  END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 99.450 0.800 99.750 ;
    END
  END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 100.050 0.800 100.350 ;
    END
  END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 100.650 0.800 100.950 ;
    END
  END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 101.250 0.800 101.550 ;
    END
  END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 101.850 0.800 102.150 ;
    END
  END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 102.450 0.800 102.750 ;
    END
  END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 103.050 0.800 103.350 ;
    END
  END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 103.650 0.800 103.950 ;
    END
  END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 104.250 0.800 104.550 ;
    END
  END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 104.850 0.800 105.150 ;
    END
  END rd_out[61]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 130.650 0.800 130.950 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 131.250 0.800 131.550 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 131.850 0.800 132.150 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 132.450 0.800 132.750 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 133.050 0.800 133.350 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 133.650 0.800 133.950 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 134.250 0.800 134.550 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 134.850 0.800 135.150 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 135.450 0.800 135.750 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 136.050 0.800 136.350 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 136.650 0.800 136.950 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 137.250 0.800 137.550 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 137.850 0.800 138.150 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 138.450 0.800 138.750 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 139.050 0.800 139.350 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 139.650 0.800 139.950 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 140.250 0.800 140.550 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 140.850 0.800 141.150 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 141.450 0.800 141.750 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 142.050 0.800 142.350 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 142.650 0.800 142.950 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 143.250 0.800 143.550 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 143.850 0.800 144.150 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 144.450 0.800 144.750 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 145.050 0.800 145.350 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 145.650 0.800 145.950 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 146.250 0.800 146.550 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 146.850 0.800 147.150 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 147.450 0.800 147.750 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 148.050 0.800 148.350 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 148.650 0.800 148.950 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 149.250 0.800 149.550 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 149.850 0.800 150.150 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 150.450 0.800 150.750 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 151.050 0.800 151.350 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 151.650 0.800 151.950 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 152.250 0.800 152.550 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 152.850 0.800 153.150 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 153.450 0.800 153.750 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 154.050 0.800 154.350 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 154.650 0.800 154.950 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 155.250 0.800 155.550 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 155.850 0.800 156.150 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 156.450 0.800 156.750 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 157.050 0.800 157.350 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 157.650 0.800 157.950 ;
    END
  END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 158.250 0.800 158.550 ;
    END
  END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 158.850 0.800 159.150 ;
    END
  END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 159.450 0.800 159.750 ;
    END
  END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 160.050 0.800 160.350 ;
    END
  END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 160.650 0.800 160.950 ;
    END
  END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 161.250 0.800 161.550 ;
    END
  END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 161.850 0.800 162.150 ;
    END
  END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 162.450 0.800 162.750 ;
    END
  END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 163.050 0.800 163.350 ;
    END
  END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 163.650 0.800 163.950 ;
    END
  END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 164.250 0.800 164.550 ;
    END
  END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 164.850 0.800 165.150 ;
    END
  END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 165.450 0.800 165.750 ;
    END
  END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 166.050 0.800 166.350 ;
    END
  END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 166.650 0.800 166.950 ;
    END
  END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 167.250 0.800 167.550 ;
    END
  END wd_in[61]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 193.050 0.800 193.350 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 193.650 0.800 193.950 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 194.250 0.800 194.550 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 194.850 0.800 195.150 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 195.450 0.800 195.750 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 196.050 0.800 196.350 ;
    END
  END addr_in[5]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 221.850 0.800 222.150 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 222.450 0.800 222.750 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 223.050 0.800 223.350 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
      RECT 5.400 6.000 6.600 227.920 ;
      RECT 15.000 6.000 16.200 227.920 ;
      RECT 24.600 6.000 25.800 227.920 ;
      RECT 34.200 6.000 35.400 227.920 ;
      RECT 43.800 6.000 45.000 227.920 ;
      RECT 53.400 6.000 54.600 227.920 ;
      RECT 63.000 6.000 64.200 227.920 ;
      RECT 72.600 6.000 73.800 227.920 ;
      RECT 82.200 6.000 83.400 227.920 ;
      RECT 91.800 6.000 93.000 227.920 ;
      RECT 101.400 6.000 102.600 227.920 ;
      RECT 111.000 6.000 112.200 227.920 ;
      RECT 120.600 6.000 121.800 227.920 ;
      RECT 130.200 6.000 131.400 227.920 ;
      RECT 139.800 6.000 141.000 227.920 ;
      RECT 149.400 6.000 150.600 227.920 ;
      RECT 159.000 6.000 160.200 227.920 ;
      RECT 168.600 6.000 169.800 227.920 ;
      RECT 178.200 6.000 179.400 227.920 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
      RECT 10.200 6.000 11.400 227.920 ;
      RECT 19.800 6.000 21.000 227.920 ;
      RECT 29.400 6.000 30.600 227.920 ;
      RECT 39.000 6.000 40.200 227.920 ;
      RECT 48.600 6.000 49.800 227.920 ;
      RECT 58.200 6.000 59.400 227.920 ;
      RECT 67.800 6.000 69.000 227.920 ;
      RECT 77.400 6.000 78.600 227.920 ;
      RECT 87.000 6.000 88.200 227.920 ;
      RECT 96.600 6.000 97.800 227.920 ;
      RECT 106.200 6.000 107.400 227.920 ;
      RECT 115.800 6.000 117.000 227.920 ;
      RECT 125.400 6.000 126.600 227.920 ;
      RECT 135.000 6.000 136.200 227.920 ;
      RECT 144.600 6.000 145.800 227.920 ;
      RECT 154.200 6.000 155.400 227.920 ;
      RECT 163.800 6.000 165.000 227.920 ;
      RECT 173.400 6.000 174.600 227.920 ;
      RECT 183.000 6.000 184.200 227.920 ;
    END
  END VDD
  OBS
    LAYER met1 ;
    RECT 0 0 189.980 233.920 ;
    LAYER met2 ;
    RECT 0 0 189.980 233.920 ;
    LAYER met3 ;
    RECT 0.800 0 189.980 233.920 ;
    RECT 0 0.000 0.800 5.850 ;
    RECT 0 6.150 0.800 6.450 ;
    RECT 0 6.750 0.800 7.050 ;
    RECT 0 7.350 0.800 7.650 ;
    RECT 0 7.950 0.800 8.250 ;
    RECT 0 8.550 0.800 8.850 ;
    RECT 0 9.150 0.800 9.450 ;
    RECT 0 9.750 0.800 10.050 ;
    RECT 0 10.350 0.800 10.650 ;
    RECT 0 10.950 0.800 11.250 ;
    RECT 0 11.550 0.800 11.850 ;
    RECT 0 12.150 0.800 12.450 ;
    RECT 0 12.750 0.800 13.050 ;
    RECT 0 13.350 0.800 13.650 ;
    RECT 0 13.950 0.800 14.250 ;
    RECT 0 14.550 0.800 14.850 ;
    RECT 0 15.150 0.800 15.450 ;
    RECT 0 15.750 0.800 16.050 ;
    RECT 0 16.350 0.800 16.650 ;
    RECT 0 16.950 0.800 17.250 ;
    RECT 0 17.550 0.800 17.850 ;
    RECT 0 18.150 0.800 18.450 ;
    RECT 0 18.750 0.800 19.050 ;
    RECT 0 19.350 0.800 19.650 ;
    RECT 0 19.950 0.800 20.250 ;
    RECT 0 20.550 0.800 20.850 ;
    RECT 0 21.150 0.800 21.450 ;
    RECT 0 21.750 0.800 22.050 ;
    RECT 0 22.350 0.800 22.650 ;
    RECT 0 22.950 0.800 23.250 ;
    RECT 0 23.550 0.800 23.850 ;
    RECT 0 24.150 0.800 24.450 ;
    RECT 0 24.750 0.800 25.050 ;
    RECT 0 25.350 0.800 25.650 ;
    RECT 0 25.950 0.800 26.250 ;
    RECT 0 26.550 0.800 26.850 ;
    RECT 0 27.150 0.800 27.450 ;
    RECT 0 27.750 0.800 28.050 ;
    RECT 0 28.350 0.800 28.650 ;
    RECT 0 28.950 0.800 29.250 ;
    RECT 0 29.550 0.800 29.850 ;
    RECT 0 30.150 0.800 30.450 ;
    RECT 0 30.750 0.800 31.050 ;
    RECT 0 31.350 0.800 31.650 ;
    RECT 0 31.950 0.800 32.250 ;
    RECT 0 32.550 0.800 32.850 ;
    RECT 0 33.150 0.800 33.450 ;
    RECT 0 33.750 0.800 34.050 ;
    RECT 0 34.350 0.800 34.650 ;
    RECT 0 34.950 0.800 35.250 ;
    RECT 0 35.550 0.800 35.850 ;
    RECT 0 36.150 0.800 36.450 ;
    RECT 0 36.750 0.800 37.050 ;
    RECT 0 37.350 0.800 37.650 ;
    RECT 0 37.950 0.800 38.250 ;
    RECT 0 38.550 0.800 38.850 ;
    RECT 0 39.150 0.800 39.450 ;
    RECT 0 39.750 0.800 40.050 ;
    RECT 0 40.350 0.800 40.650 ;
    RECT 0 40.950 0.800 41.250 ;
    RECT 0 41.550 0.800 41.850 ;
    RECT 0 42.150 0.800 42.450 ;
    RECT 0 42.750 0.800 68.250 ;
    RECT 0 68.550 0.800 68.850 ;
    RECT 0 69.150 0.800 69.450 ;
    RECT 0 69.750 0.800 70.050 ;
    RECT 0 70.350 0.800 70.650 ;
    RECT 0 70.950 0.800 71.250 ;
    RECT 0 71.550 0.800 71.850 ;
    RECT 0 72.150 0.800 72.450 ;
    RECT 0 72.750 0.800 73.050 ;
    RECT 0 73.350 0.800 73.650 ;
    RECT 0 73.950 0.800 74.250 ;
    RECT 0 74.550 0.800 74.850 ;
    RECT 0 75.150 0.800 75.450 ;
    RECT 0 75.750 0.800 76.050 ;
    RECT 0 76.350 0.800 76.650 ;
    RECT 0 76.950 0.800 77.250 ;
    RECT 0 77.550 0.800 77.850 ;
    RECT 0 78.150 0.800 78.450 ;
    RECT 0 78.750 0.800 79.050 ;
    RECT 0 79.350 0.800 79.650 ;
    RECT 0 79.950 0.800 80.250 ;
    RECT 0 80.550 0.800 80.850 ;
    RECT 0 81.150 0.800 81.450 ;
    RECT 0 81.750 0.800 82.050 ;
    RECT 0 82.350 0.800 82.650 ;
    RECT 0 82.950 0.800 83.250 ;
    RECT 0 83.550 0.800 83.850 ;
    RECT 0 84.150 0.800 84.450 ;
    RECT 0 84.750 0.800 85.050 ;
    RECT 0 85.350 0.800 85.650 ;
    RECT 0 85.950 0.800 86.250 ;
    RECT 0 86.550 0.800 86.850 ;
    RECT 0 87.150 0.800 87.450 ;
    RECT 0 87.750 0.800 88.050 ;
    RECT 0 88.350 0.800 88.650 ;
    RECT 0 88.950 0.800 89.250 ;
    RECT 0 89.550 0.800 89.850 ;
    RECT 0 90.150 0.800 90.450 ;
    RECT 0 90.750 0.800 91.050 ;
    RECT 0 91.350 0.800 91.650 ;
    RECT 0 91.950 0.800 92.250 ;
    RECT 0 92.550 0.800 92.850 ;
    RECT 0 93.150 0.800 93.450 ;
    RECT 0 93.750 0.800 94.050 ;
    RECT 0 94.350 0.800 94.650 ;
    RECT 0 94.950 0.800 95.250 ;
    RECT 0 95.550 0.800 95.850 ;
    RECT 0 96.150 0.800 96.450 ;
    RECT 0 96.750 0.800 97.050 ;
    RECT 0 97.350 0.800 97.650 ;
    RECT 0 97.950 0.800 98.250 ;
    RECT 0 98.550 0.800 98.850 ;
    RECT 0 99.150 0.800 99.450 ;
    RECT 0 99.750 0.800 100.050 ;
    RECT 0 100.350 0.800 100.650 ;
    RECT 0 100.950 0.800 101.250 ;
    RECT 0 101.550 0.800 101.850 ;
    RECT 0 102.150 0.800 102.450 ;
    RECT 0 102.750 0.800 103.050 ;
    RECT 0 103.350 0.800 103.650 ;
    RECT 0 103.950 0.800 104.250 ;
    RECT 0 104.550 0.800 104.850 ;
    RECT 0 105.150 0.800 130.650 ;
    RECT 0 130.950 0.800 131.250 ;
    RECT 0 131.550 0.800 131.850 ;
    RECT 0 132.150 0.800 132.450 ;
    RECT 0 132.750 0.800 133.050 ;
    RECT 0 133.350 0.800 133.650 ;
    RECT 0 133.950 0.800 134.250 ;
    RECT 0 134.550 0.800 134.850 ;
    RECT 0 135.150 0.800 135.450 ;
    RECT 0 135.750 0.800 136.050 ;
    RECT 0 136.350 0.800 136.650 ;
    RECT 0 136.950 0.800 137.250 ;
    RECT 0 137.550 0.800 137.850 ;
    RECT 0 138.150 0.800 138.450 ;
    RECT 0 138.750 0.800 139.050 ;
    RECT 0 139.350 0.800 139.650 ;
    RECT 0 139.950 0.800 140.250 ;
    RECT 0 140.550 0.800 140.850 ;
    RECT 0 141.150 0.800 141.450 ;
    RECT 0 141.750 0.800 142.050 ;
    RECT 0 142.350 0.800 142.650 ;
    RECT 0 142.950 0.800 143.250 ;
    RECT 0 143.550 0.800 143.850 ;
    RECT 0 144.150 0.800 144.450 ;
    RECT 0 144.750 0.800 145.050 ;
    RECT 0 145.350 0.800 145.650 ;
    RECT 0 145.950 0.800 146.250 ;
    RECT 0 146.550 0.800 146.850 ;
    RECT 0 147.150 0.800 147.450 ;
    RECT 0 147.750 0.800 148.050 ;
    RECT 0 148.350 0.800 148.650 ;
    RECT 0 148.950 0.800 149.250 ;
    RECT 0 149.550 0.800 149.850 ;
    RECT 0 150.150 0.800 150.450 ;
    RECT 0 150.750 0.800 151.050 ;
    RECT 0 151.350 0.800 151.650 ;
    RECT 0 151.950 0.800 152.250 ;
    RECT 0 152.550 0.800 152.850 ;
    RECT 0 153.150 0.800 153.450 ;
    RECT 0 153.750 0.800 154.050 ;
    RECT 0 154.350 0.800 154.650 ;
    RECT 0 154.950 0.800 155.250 ;
    RECT 0 155.550 0.800 155.850 ;
    RECT 0 156.150 0.800 156.450 ;
    RECT 0 156.750 0.800 157.050 ;
    RECT 0 157.350 0.800 157.650 ;
    RECT 0 157.950 0.800 158.250 ;
    RECT 0 158.550 0.800 158.850 ;
    RECT 0 159.150 0.800 159.450 ;
    RECT 0 159.750 0.800 160.050 ;
    RECT 0 160.350 0.800 160.650 ;
    RECT 0 160.950 0.800 161.250 ;
    RECT 0 161.550 0.800 161.850 ;
    RECT 0 162.150 0.800 162.450 ;
    RECT 0 162.750 0.800 163.050 ;
    RECT 0 163.350 0.800 163.650 ;
    RECT 0 163.950 0.800 164.250 ;
    RECT 0 164.550 0.800 164.850 ;
    RECT 0 165.150 0.800 165.450 ;
    RECT 0 165.750 0.800 166.050 ;
    RECT 0 166.350 0.800 166.650 ;
    RECT 0 166.950 0.800 167.250 ;
    RECT 0 167.550 0.800 193.050 ;
    RECT 0 193.350 0.800 193.650 ;
    RECT 0 193.950 0.800 194.250 ;
    RECT 0 194.550 0.800 194.850 ;
    RECT 0 195.150 0.800 195.450 ;
    RECT 0 195.750 0.800 196.050 ;
    RECT 0 196.350 0.800 221.850 ;
    RECT 0 222.150 0.800 222.450 ;
    RECT 0 222.750 0.800 223.050 ;
    RECT 0 223.350 0.800 233.920 ;
    LAYER met4 ;
    RECT 0 0 189.980 6.000 ;
    RECT 0 227.920 189.980 233.920 ;
    RECT 0.000 6.000 5.400 227.920 ;
    RECT 6.600 6.000 10.200 227.920 ;
    RECT 11.400 6.000 15.000 227.920 ;
    RECT 16.200 6.000 19.800 227.920 ;
    RECT 21.000 6.000 24.600 227.920 ;
    RECT 25.800 6.000 29.400 227.920 ;
    RECT 30.600 6.000 34.200 227.920 ;
    RECT 35.400 6.000 39.000 227.920 ;
    RECT 40.200 6.000 43.800 227.920 ;
    RECT 45.000 6.000 48.600 227.920 ;
    RECT 49.800 6.000 53.400 227.920 ;
    RECT 54.600 6.000 58.200 227.920 ;
    RECT 59.400 6.000 63.000 227.920 ;
    RECT 64.200 6.000 67.800 227.920 ;
    RECT 69.000 6.000 72.600 227.920 ;
    RECT 73.800 6.000 77.400 227.920 ;
    RECT 78.600 6.000 82.200 227.920 ;
    RECT 83.400 6.000 87.000 227.920 ;
    RECT 88.200 6.000 91.800 227.920 ;
    RECT 93.000 6.000 96.600 227.920 ;
    RECT 97.800 6.000 101.400 227.920 ;
    RECT 102.600 6.000 106.200 227.920 ;
    RECT 107.400 6.000 111.000 227.920 ;
    RECT 112.200 6.000 115.800 227.920 ;
    RECT 117.000 6.000 120.600 227.920 ;
    RECT 121.800 6.000 125.400 227.920 ;
    RECT 126.600 6.000 130.200 227.920 ;
    RECT 131.400 6.000 135.000 227.920 ;
    RECT 136.200 6.000 139.800 227.920 ;
    RECT 141.000 6.000 144.600 227.920 ;
    RECT 145.800 6.000 149.400 227.920 ;
    RECT 150.600 6.000 154.200 227.920 ;
    RECT 155.400 6.000 159.000 227.920 ;
    RECT 160.200 6.000 163.800 227.920 ;
    RECT 165.000 6.000 168.600 227.920 ;
    RECT 169.800 6.000 173.400 227.920 ;
    RECT 174.600 6.000 178.200 227.920 ;
    RECT 179.400 6.000 183.000 227.920 ;
    RECT 184.200 6.000 189.980 227.920 ;
    LAYER OVERLAP ;
    RECT 0 0 189.980 233.920 ;
  END
END fakeram130_64x62

END LIBRARY
