VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram130_1024x32
  FOREIGN fakeram130_1024x32 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 540.040 BY 440.640 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 5.850 0.800 6.150 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 9.450 0.800 9.750 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 13.050 0.800 13.350 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 16.650 0.800 16.950 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 20.250 0.800 20.550 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 23.850 0.800 24.150 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 27.450 0.800 27.750 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 31.050 0.800 31.350 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 34.650 0.800 34.950 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 38.250 0.800 38.550 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 41.850 0.800 42.150 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 45.450 0.800 45.750 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 49.050 0.800 49.350 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 52.650 0.800 52.950 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 56.250 0.800 56.550 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 59.850 0.800 60.150 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 63.450 0.800 63.750 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 67.050 0.800 67.350 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 70.650 0.800 70.950 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 74.250 0.800 74.550 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 77.850 0.800 78.150 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 81.450 0.800 81.750 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 85.050 0.800 85.350 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 88.650 0.800 88.950 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 92.250 0.800 92.550 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 95.850 0.800 96.150 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 99.450 0.800 99.750 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 103.050 0.800 103.350 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 106.650 0.800 106.950 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 110.250 0.800 110.550 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 113.850 0.800 114.150 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 117.450 0.800 117.750 ;
    END
  END w_mask_in[31]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 126.450 0.800 126.750 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 130.050 0.800 130.350 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 133.650 0.800 133.950 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 137.250 0.800 137.550 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 140.850 0.800 141.150 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 144.450 0.800 144.750 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 148.050 0.800 148.350 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 151.650 0.800 151.950 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 155.250 0.800 155.550 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 158.850 0.800 159.150 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 162.450 0.800 162.750 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 166.050 0.800 166.350 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 169.650 0.800 169.950 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 173.250 0.800 173.550 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 176.850 0.800 177.150 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 180.450 0.800 180.750 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 184.050 0.800 184.350 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 187.650 0.800 187.950 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 191.250 0.800 191.550 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 194.850 0.800 195.150 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 198.450 0.800 198.750 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 202.050 0.800 202.350 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 205.650 0.800 205.950 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 209.250 0.800 209.550 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 212.850 0.800 213.150 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 216.450 0.800 216.750 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 220.050 0.800 220.350 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 223.650 0.800 223.950 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 227.250 0.800 227.550 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 230.850 0.800 231.150 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 234.450 0.800 234.750 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 238.050 0.800 238.350 ;
    END
  END rd_out[31]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 247.050 0.800 247.350 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 250.650 0.800 250.950 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 254.250 0.800 254.550 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 257.850 0.800 258.150 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 261.450 0.800 261.750 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 265.050 0.800 265.350 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 268.650 0.800 268.950 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 272.250 0.800 272.550 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 275.850 0.800 276.150 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 279.450 0.800 279.750 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 283.050 0.800 283.350 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 286.650 0.800 286.950 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 290.250 0.800 290.550 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 293.850 0.800 294.150 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 297.450 0.800 297.750 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 301.050 0.800 301.350 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 304.650 0.800 304.950 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 308.250 0.800 308.550 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 311.850 0.800 312.150 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 315.450 0.800 315.750 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 319.050 0.800 319.350 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 322.650 0.800 322.950 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 326.250 0.800 326.550 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 329.850 0.800 330.150 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 333.450 0.800 333.750 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 337.050 0.800 337.350 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 340.650 0.800 340.950 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 344.250 0.800 344.550 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 347.850 0.800 348.150 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 351.450 0.800 351.750 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 355.050 0.800 355.350 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 358.650 0.800 358.950 ;
    END
  END wd_in[31]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 367.650 0.800 367.950 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 371.250 0.800 371.550 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 374.850 0.800 375.150 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 378.450 0.800 378.750 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 382.050 0.800 382.350 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 385.650 0.800 385.950 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 389.250 0.800 389.550 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 392.850 0.800 393.150 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 396.450 0.800 396.750 ;
    END
  END addr_in[8]
  PIN addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 400.050 0.800 400.350 ;
    END
  END addr_in[9]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 409.050 0.800 409.350 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 412.650 0.800 412.950 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 416.250 0.800 416.550 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
      RECT 5.400 6.000 6.600 434.640 ;
      RECT 15.000 6.000 16.200 434.640 ;
      RECT 24.600 6.000 25.800 434.640 ;
      RECT 34.200 6.000 35.400 434.640 ;
      RECT 43.800 6.000 45.000 434.640 ;
      RECT 53.400 6.000 54.600 434.640 ;
      RECT 63.000 6.000 64.200 434.640 ;
      RECT 72.600 6.000 73.800 434.640 ;
      RECT 82.200 6.000 83.400 434.640 ;
      RECT 91.800 6.000 93.000 434.640 ;
      RECT 101.400 6.000 102.600 434.640 ;
      RECT 111.000 6.000 112.200 434.640 ;
      RECT 120.600 6.000 121.800 434.640 ;
      RECT 130.200 6.000 131.400 434.640 ;
      RECT 139.800 6.000 141.000 434.640 ;
      RECT 149.400 6.000 150.600 434.640 ;
      RECT 159.000 6.000 160.200 434.640 ;
      RECT 168.600 6.000 169.800 434.640 ;
      RECT 178.200 6.000 179.400 434.640 ;
      RECT 187.800 6.000 189.000 434.640 ;
      RECT 197.400 6.000 198.600 434.640 ;
      RECT 207.000 6.000 208.200 434.640 ;
      RECT 216.600 6.000 217.800 434.640 ;
      RECT 226.200 6.000 227.400 434.640 ;
      RECT 235.800 6.000 237.000 434.640 ;
      RECT 245.400 6.000 246.600 434.640 ;
      RECT 255.000 6.000 256.200 434.640 ;
      RECT 264.600 6.000 265.800 434.640 ;
      RECT 274.200 6.000 275.400 434.640 ;
      RECT 283.800 6.000 285.000 434.640 ;
      RECT 293.400 6.000 294.600 434.640 ;
      RECT 303.000 6.000 304.200 434.640 ;
      RECT 312.600 6.000 313.800 434.640 ;
      RECT 322.200 6.000 323.400 434.640 ;
      RECT 331.800 6.000 333.000 434.640 ;
      RECT 341.400 6.000 342.600 434.640 ;
      RECT 351.000 6.000 352.200 434.640 ;
      RECT 360.600 6.000 361.800 434.640 ;
      RECT 370.200 6.000 371.400 434.640 ;
      RECT 379.800 6.000 381.000 434.640 ;
      RECT 389.400 6.000 390.600 434.640 ;
      RECT 399.000 6.000 400.200 434.640 ;
      RECT 408.600 6.000 409.800 434.640 ;
      RECT 418.200 6.000 419.400 434.640 ;
      RECT 427.800 6.000 429.000 434.640 ;
      RECT 437.400 6.000 438.600 434.640 ;
      RECT 447.000 6.000 448.200 434.640 ;
      RECT 456.600 6.000 457.800 434.640 ;
      RECT 466.200 6.000 467.400 434.640 ;
      RECT 475.800 6.000 477.000 434.640 ;
      RECT 485.400 6.000 486.600 434.640 ;
      RECT 495.000 6.000 496.200 434.640 ;
      RECT 504.600 6.000 505.800 434.640 ;
      RECT 514.200 6.000 515.400 434.640 ;
      RECT 523.800 6.000 525.000 434.640 ;
      RECT 533.400 6.000 534.600 434.640 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
      RECT 10.200 6.000 11.400 434.640 ;
      RECT 19.800 6.000 21.000 434.640 ;
      RECT 29.400 6.000 30.600 434.640 ;
      RECT 39.000 6.000 40.200 434.640 ;
      RECT 48.600 6.000 49.800 434.640 ;
      RECT 58.200 6.000 59.400 434.640 ;
      RECT 67.800 6.000 69.000 434.640 ;
      RECT 77.400 6.000 78.600 434.640 ;
      RECT 87.000 6.000 88.200 434.640 ;
      RECT 96.600 6.000 97.800 434.640 ;
      RECT 106.200 6.000 107.400 434.640 ;
      RECT 115.800 6.000 117.000 434.640 ;
      RECT 125.400 6.000 126.600 434.640 ;
      RECT 135.000 6.000 136.200 434.640 ;
      RECT 144.600 6.000 145.800 434.640 ;
      RECT 154.200 6.000 155.400 434.640 ;
      RECT 163.800 6.000 165.000 434.640 ;
      RECT 173.400 6.000 174.600 434.640 ;
      RECT 183.000 6.000 184.200 434.640 ;
      RECT 192.600 6.000 193.800 434.640 ;
      RECT 202.200 6.000 203.400 434.640 ;
      RECT 211.800 6.000 213.000 434.640 ;
      RECT 221.400 6.000 222.600 434.640 ;
      RECT 231.000 6.000 232.200 434.640 ;
      RECT 240.600 6.000 241.800 434.640 ;
      RECT 250.200 6.000 251.400 434.640 ;
      RECT 259.800 6.000 261.000 434.640 ;
      RECT 269.400 6.000 270.600 434.640 ;
      RECT 279.000 6.000 280.200 434.640 ;
      RECT 288.600 6.000 289.800 434.640 ;
      RECT 298.200 6.000 299.400 434.640 ;
      RECT 307.800 6.000 309.000 434.640 ;
      RECT 317.400 6.000 318.600 434.640 ;
      RECT 327.000 6.000 328.200 434.640 ;
      RECT 336.600 6.000 337.800 434.640 ;
      RECT 346.200 6.000 347.400 434.640 ;
      RECT 355.800 6.000 357.000 434.640 ;
      RECT 365.400 6.000 366.600 434.640 ;
      RECT 375.000 6.000 376.200 434.640 ;
      RECT 384.600 6.000 385.800 434.640 ;
      RECT 394.200 6.000 395.400 434.640 ;
      RECT 403.800 6.000 405.000 434.640 ;
      RECT 413.400 6.000 414.600 434.640 ;
      RECT 423.000 6.000 424.200 434.640 ;
      RECT 432.600 6.000 433.800 434.640 ;
      RECT 442.200 6.000 443.400 434.640 ;
      RECT 451.800 6.000 453.000 434.640 ;
      RECT 461.400 6.000 462.600 434.640 ;
      RECT 471.000 6.000 472.200 434.640 ;
      RECT 480.600 6.000 481.800 434.640 ;
      RECT 490.200 6.000 491.400 434.640 ;
      RECT 499.800 6.000 501.000 434.640 ;
      RECT 509.400 6.000 510.600 434.640 ;
      RECT 519.000 6.000 520.200 434.640 ;
      RECT 528.600 6.000 529.800 434.640 ;
    END
  END VDD
  OBS
    LAYER met1 ;
    RECT 0 0 540.040 440.640 ;
    LAYER met2 ;
    RECT 0 0 540.040 440.640 ;
    LAYER met3 ;
    RECT 0.800 0 540.040 440.640 ;
    RECT 0 0.000 0.800 5.850 ;
    RECT 0 6.150 0.800 9.450 ;
    RECT 0 9.750 0.800 13.050 ;
    RECT 0 13.350 0.800 16.650 ;
    RECT 0 16.950 0.800 20.250 ;
    RECT 0 20.550 0.800 23.850 ;
    RECT 0 24.150 0.800 27.450 ;
    RECT 0 27.750 0.800 31.050 ;
    RECT 0 31.350 0.800 34.650 ;
    RECT 0 34.950 0.800 38.250 ;
    RECT 0 38.550 0.800 41.850 ;
    RECT 0 42.150 0.800 45.450 ;
    RECT 0 45.750 0.800 49.050 ;
    RECT 0 49.350 0.800 52.650 ;
    RECT 0 52.950 0.800 56.250 ;
    RECT 0 56.550 0.800 59.850 ;
    RECT 0 60.150 0.800 63.450 ;
    RECT 0 63.750 0.800 67.050 ;
    RECT 0 67.350 0.800 70.650 ;
    RECT 0 70.950 0.800 74.250 ;
    RECT 0 74.550 0.800 77.850 ;
    RECT 0 78.150 0.800 81.450 ;
    RECT 0 81.750 0.800 85.050 ;
    RECT 0 85.350 0.800 88.650 ;
    RECT 0 88.950 0.800 92.250 ;
    RECT 0 92.550 0.800 95.850 ;
    RECT 0 96.150 0.800 99.450 ;
    RECT 0 99.750 0.800 103.050 ;
    RECT 0 103.350 0.800 106.650 ;
    RECT 0 106.950 0.800 110.250 ;
    RECT 0 110.550 0.800 113.850 ;
    RECT 0 114.150 0.800 117.450 ;
    RECT 0 117.750 0.800 126.450 ;
    RECT 0 126.750 0.800 130.050 ;
    RECT 0 130.350 0.800 133.650 ;
    RECT 0 133.950 0.800 137.250 ;
    RECT 0 137.550 0.800 140.850 ;
    RECT 0 141.150 0.800 144.450 ;
    RECT 0 144.750 0.800 148.050 ;
    RECT 0 148.350 0.800 151.650 ;
    RECT 0 151.950 0.800 155.250 ;
    RECT 0 155.550 0.800 158.850 ;
    RECT 0 159.150 0.800 162.450 ;
    RECT 0 162.750 0.800 166.050 ;
    RECT 0 166.350 0.800 169.650 ;
    RECT 0 169.950 0.800 173.250 ;
    RECT 0 173.550 0.800 176.850 ;
    RECT 0 177.150 0.800 180.450 ;
    RECT 0 180.750 0.800 184.050 ;
    RECT 0 184.350 0.800 187.650 ;
    RECT 0 187.950 0.800 191.250 ;
    RECT 0 191.550 0.800 194.850 ;
    RECT 0 195.150 0.800 198.450 ;
    RECT 0 198.750 0.800 202.050 ;
    RECT 0 202.350 0.800 205.650 ;
    RECT 0 205.950 0.800 209.250 ;
    RECT 0 209.550 0.800 212.850 ;
    RECT 0 213.150 0.800 216.450 ;
    RECT 0 216.750 0.800 220.050 ;
    RECT 0 220.350 0.800 223.650 ;
    RECT 0 223.950 0.800 227.250 ;
    RECT 0 227.550 0.800 230.850 ;
    RECT 0 231.150 0.800 234.450 ;
    RECT 0 234.750 0.800 238.050 ;
    RECT 0 238.350 0.800 247.050 ;
    RECT 0 247.350 0.800 250.650 ;
    RECT 0 250.950 0.800 254.250 ;
    RECT 0 254.550 0.800 257.850 ;
    RECT 0 258.150 0.800 261.450 ;
    RECT 0 261.750 0.800 265.050 ;
    RECT 0 265.350 0.800 268.650 ;
    RECT 0 268.950 0.800 272.250 ;
    RECT 0 272.550 0.800 275.850 ;
    RECT 0 276.150 0.800 279.450 ;
    RECT 0 279.750 0.800 283.050 ;
    RECT 0 283.350 0.800 286.650 ;
    RECT 0 286.950 0.800 290.250 ;
    RECT 0 290.550 0.800 293.850 ;
    RECT 0 294.150 0.800 297.450 ;
    RECT 0 297.750 0.800 301.050 ;
    RECT 0 301.350 0.800 304.650 ;
    RECT 0 304.950 0.800 308.250 ;
    RECT 0 308.550 0.800 311.850 ;
    RECT 0 312.150 0.800 315.450 ;
    RECT 0 315.750 0.800 319.050 ;
    RECT 0 319.350 0.800 322.650 ;
    RECT 0 322.950 0.800 326.250 ;
    RECT 0 326.550 0.800 329.850 ;
    RECT 0 330.150 0.800 333.450 ;
    RECT 0 333.750 0.800 337.050 ;
    RECT 0 337.350 0.800 340.650 ;
    RECT 0 340.950 0.800 344.250 ;
    RECT 0 344.550 0.800 347.850 ;
    RECT 0 348.150 0.800 351.450 ;
    RECT 0 351.750 0.800 355.050 ;
    RECT 0 355.350 0.800 358.650 ;
    RECT 0 358.950 0.800 367.650 ;
    RECT 0 367.950 0.800 371.250 ;
    RECT 0 371.550 0.800 374.850 ;
    RECT 0 375.150 0.800 378.450 ;
    RECT 0 378.750 0.800 382.050 ;
    RECT 0 382.350 0.800 385.650 ;
    RECT 0 385.950 0.800 389.250 ;
    RECT 0 389.550 0.800 392.850 ;
    RECT 0 393.150 0.800 396.450 ;
    RECT 0 396.750 0.800 400.050 ;
    RECT 0 400.350 0.800 409.050 ;
    RECT 0 409.350 0.800 412.650 ;
    RECT 0 412.950 0.800 416.250 ;
    RECT 0 416.550 0.800 440.640 ;
    LAYER met4 ;
    RECT 0 0 540.040 6.000 ;
    RECT 0 434.640 540.040 440.640 ;
    RECT 0.000 6.000 5.400 434.640 ;
    RECT 6.600 6.000 10.200 434.640 ;
    RECT 11.400 6.000 15.000 434.640 ;
    RECT 16.200 6.000 19.800 434.640 ;
    RECT 21.000 6.000 24.600 434.640 ;
    RECT 25.800 6.000 29.400 434.640 ;
    RECT 30.600 6.000 34.200 434.640 ;
    RECT 35.400 6.000 39.000 434.640 ;
    RECT 40.200 6.000 43.800 434.640 ;
    RECT 45.000 6.000 48.600 434.640 ;
    RECT 49.800 6.000 53.400 434.640 ;
    RECT 54.600 6.000 58.200 434.640 ;
    RECT 59.400 6.000 63.000 434.640 ;
    RECT 64.200 6.000 67.800 434.640 ;
    RECT 69.000 6.000 72.600 434.640 ;
    RECT 73.800 6.000 77.400 434.640 ;
    RECT 78.600 6.000 82.200 434.640 ;
    RECT 83.400 6.000 87.000 434.640 ;
    RECT 88.200 6.000 91.800 434.640 ;
    RECT 93.000 6.000 96.600 434.640 ;
    RECT 97.800 6.000 101.400 434.640 ;
    RECT 102.600 6.000 106.200 434.640 ;
    RECT 107.400 6.000 111.000 434.640 ;
    RECT 112.200 6.000 115.800 434.640 ;
    RECT 117.000 6.000 120.600 434.640 ;
    RECT 121.800 6.000 125.400 434.640 ;
    RECT 126.600 6.000 130.200 434.640 ;
    RECT 131.400 6.000 135.000 434.640 ;
    RECT 136.200 6.000 139.800 434.640 ;
    RECT 141.000 6.000 144.600 434.640 ;
    RECT 145.800 6.000 149.400 434.640 ;
    RECT 150.600 6.000 154.200 434.640 ;
    RECT 155.400 6.000 159.000 434.640 ;
    RECT 160.200 6.000 163.800 434.640 ;
    RECT 165.000 6.000 168.600 434.640 ;
    RECT 169.800 6.000 173.400 434.640 ;
    RECT 174.600 6.000 178.200 434.640 ;
    RECT 179.400 6.000 183.000 434.640 ;
    RECT 184.200 6.000 187.800 434.640 ;
    RECT 189.000 6.000 192.600 434.640 ;
    RECT 193.800 6.000 197.400 434.640 ;
    RECT 198.600 6.000 202.200 434.640 ;
    RECT 203.400 6.000 207.000 434.640 ;
    RECT 208.200 6.000 211.800 434.640 ;
    RECT 213.000 6.000 216.600 434.640 ;
    RECT 217.800 6.000 221.400 434.640 ;
    RECT 222.600 6.000 226.200 434.640 ;
    RECT 227.400 6.000 231.000 434.640 ;
    RECT 232.200 6.000 235.800 434.640 ;
    RECT 237.000 6.000 240.600 434.640 ;
    RECT 241.800 6.000 245.400 434.640 ;
    RECT 246.600 6.000 250.200 434.640 ;
    RECT 251.400 6.000 255.000 434.640 ;
    RECT 256.200 6.000 259.800 434.640 ;
    RECT 261.000 6.000 264.600 434.640 ;
    RECT 265.800 6.000 269.400 434.640 ;
    RECT 270.600 6.000 274.200 434.640 ;
    RECT 275.400 6.000 279.000 434.640 ;
    RECT 280.200 6.000 283.800 434.640 ;
    RECT 285.000 6.000 288.600 434.640 ;
    RECT 289.800 6.000 293.400 434.640 ;
    RECT 294.600 6.000 298.200 434.640 ;
    RECT 299.400 6.000 303.000 434.640 ;
    RECT 304.200 6.000 307.800 434.640 ;
    RECT 309.000 6.000 312.600 434.640 ;
    RECT 313.800 6.000 317.400 434.640 ;
    RECT 318.600 6.000 322.200 434.640 ;
    RECT 323.400 6.000 327.000 434.640 ;
    RECT 328.200 6.000 331.800 434.640 ;
    RECT 333.000 6.000 336.600 434.640 ;
    RECT 337.800 6.000 341.400 434.640 ;
    RECT 342.600 6.000 346.200 434.640 ;
    RECT 347.400 6.000 351.000 434.640 ;
    RECT 352.200 6.000 355.800 434.640 ;
    RECT 357.000 6.000 360.600 434.640 ;
    RECT 361.800 6.000 365.400 434.640 ;
    RECT 366.600 6.000 370.200 434.640 ;
    RECT 371.400 6.000 375.000 434.640 ;
    RECT 376.200 6.000 379.800 434.640 ;
    RECT 381.000 6.000 384.600 434.640 ;
    RECT 385.800 6.000 389.400 434.640 ;
    RECT 390.600 6.000 394.200 434.640 ;
    RECT 395.400 6.000 399.000 434.640 ;
    RECT 400.200 6.000 403.800 434.640 ;
    RECT 405.000 6.000 408.600 434.640 ;
    RECT 409.800 6.000 413.400 434.640 ;
    RECT 414.600 6.000 418.200 434.640 ;
    RECT 419.400 6.000 423.000 434.640 ;
    RECT 424.200 6.000 427.800 434.640 ;
    RECT 429.000 6.000 432.600 434.640 ;
    RECT 433.800 6.000 437.400 434.640 ;
    RECT 438.600 6.000 442.200 434.640 ;
    RECT 443.400 6.000 447.000 434.640 ;
    RECT 448.200 6.000 451.800 434.640 ;
    RECT 453.000 6.000 456.600 434.640 ;
    RECT 457.800 6.000 461.400 434.640 ;
    RECT 462.600 6.000 466.200 434.640 ;
    RECT 467.400 6.000 471.000 434.640 ;
    RECT 472.200 6.000 475.800 434.640 ;
    RECT 477.000 6.000 480.600 434.640 ;
    RECT 481.800 6.000 485.400 434.640 ;
    RECT 486.600 6.000 490.200 434.640 ;
    RECT 491.400 6.000 495.000 434.640 ;
    RECT 496.200 6.000 499.800 434.640 ;
    RECT 501.000 6.000 504.600 434.640 ;
    RECT 505.800 6.000 509.400 434.640 ;
    RECT 510.600 6.000 514.200 434.640 ;
    RECT 515.400 6.000 519.000 434.640 ;
    RECT 520.200 6.000 523.800 434.640 ;
    RECT 525.000 6.000 528.600 434.640 ;
    RECT 529.800 6.000 533.400 434.640 ;
    RECT 534.600 6.000 540.040 434.640 ;
    LAYER OVERLAP ;
    RECT 0 0 540.040 440.640 ;
  END
END fakeram130_1024x32

END LIBRARY
