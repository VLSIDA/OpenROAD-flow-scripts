VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram130_64x15
  FOREIGN fakeram130_64x15 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 281.060 BY 73.440 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 5.850 0.800 6.150 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 6.450 0.800 6.750 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 7.050 0.800 7.350 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 7.650 0.800 7.950 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 8.250 0.800 8.550 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 8.850 0.800 9.150 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 9.450 0.800 9.750 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 10.050 0.800 10.350 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 10.650 0.800 10.950 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 11.250 0.800 11.550 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 11.850 0.800 12.150 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 12.450 0.800 12.750 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 13.050 0.800 13.350 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 13.650 0.800 13.950 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 14.250 0.800 14.550 ;
    END
  END w_mask_in[14]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 21.450 0.800 21.750 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 22.050 0.800 22.350 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 22.650 0.800 22.950 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 23.250 0.800 23.550 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 23.850 0.800 24.150 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 24.450 0.800 24.750 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 25.050 0.800 25.350 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 25.650 0.800 25.950 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 26.250 0.800 26.550 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 26.850 0.800 27.150 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 27.450 0.800 27.750 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 28.050 0.800 28.350 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 28.650 0.800 28.950 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 29.250 0.800 29.550 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 29.850 0.800 30.150 ;
    END
  END rd_out[14]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 37.050 0.800 37.350 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 37.650 0.800 37.950 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 38.250 0.800 38.550 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 38.850 0.800 39.150 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 39.450 0.800 39.750 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 40.050 0.800 40.350 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 40.650 0.800 40.950 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 41.250 0.800 41.550 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 41.850 0.800 42.150 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 42.450 0.800 42.750 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 43.050 0.800 43.350 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 43.650 0.800 43.950 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 44.250 0.800 44.550 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 44.850 0.800 45.150 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 45.450 0.800 45.750 ;
    END
  END wd_in[14]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 52.650 0.800 52.950 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 53.250 0.800 53.550 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 53.850 0.800 54.150 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 54.450 0.800 54.750 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 55.050 0.800 55.350 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 55.650 0.800 55.950 ;
    END
  END addr_in[5]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 62.850 0.800 63.150 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 63.450 0.800 63.750 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 64.050 0.800 64.350 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
      RECT 5.400 6.000 6.600 67.440 ;
      RECT 15.000 6.000 16.200 67.440 ;
      RECT 24.600 6.000 25.800 67.440 ;
      RECT 34.200 6.000 35.400 67.440 ;
      RECT 43.800 6.000 45.000 67.440 ;
      RECT 53.400 6.000 54.600 67.440 ;
      RECT 63.000 6.000 64.200 67.440 ;
      RECT 72.600 6.000 73.800 67.440 ;
      RECT 82.200 6.000 83.400 67.440 ;
      RECT 91.800 6.000 93.000 67.440 ;
      RECT 101.400 6.000 102.600 67.440 ;
      RECT 111.000 6.000 112.200 67.440 ;
      RECT 120.600 6.000 121.800 67.440 ;
      RECT 130.200 6.000 131.400 67.440 ;
      RECT 139.800 6.000 141.000 67.440 ;
      RECT 149.400 6.000 150.600 67.440 ;
      RECT 159.000 6.000 160.200 67.440 ;
      RECT 168.600 6.000 169.800 67.440 ;
      RECT 178.200 6.000 179.400 67.440 ;
      RECT 187.800 6.000 189.000 67.440 ;
      RECT 197.400 6.000 198.600 67.440 ;
      RECT 207.000 6.000 208.200 67.440 ;
      RECT 216.600 6.000 217.800 67.440 ;
      RECT 226.200 6.000 227.400 67.440 ;
      RECT 235.800 6.000 237.000 67.440 ;
      RECT 245.400 6.000 246.600 67.440 ;
      RECT 255.000 6.000 256.200 67.440 ;
      RECT 264.600 6.000 265.800 67.440 ;
      RECT 274.200 6.000 275.400 67.440 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
      RECT 10.200 6.000 11.400 67.440 ;
      RECT 19.800 6.000 21.000 67.440 ;
      RECT 29.400 6.000 30.600 67.440 ;
      RECT 39.000 6.000 40.200 67.440 ;
      RECT 48.600 6.000 49.800 67.440 ;
      RECT 58.200 6.000 59.400 67.440 ;
      RECT 67.800 6.000 69.000 67.440 ;
      RECT 77.400 6.000 78.600 67.440 ;
      RECT 87.000 6.000 88.200 67.440 ;
      RECT 96.600 6.000 97.800 67.440 ;
      RECT 106.200 6.000 107.400 67.440 ;
      RECT 115.800 6.000 117.000 67.440 ;
      RECT 125.400 6.000 126.600 67.440 ;
      RECT 135.000 6.000 136.200 67.440 ;
      RECT 144.600 6.000 145.800 67.440 ;
      RECT 154.200 6.000 155.400 67.440 ;
      RECT 163.800 6.000 165.000 67.440 ;
      RECT 173.400 6.000 174.600 67.440 ;
      RECT 183.000 6.000 184.200 67.440 ;
      RECT 192.600 6.000 193.800 67.440 ;
      RECT 202.200 6.000 203.400 67.440 ;
      RECT 211.800 6.000 213.000 67.440 ;
      RECT 221.400 6.000 222.600 67.440 ;
      RECT 231.000 6.000 232.200 67.440 ;
      RECT 240.600 6.000 241.800 67.440 ;
      RECT 250.200 6.000 251.400 67.440 ;
      RECT 259.800 6.000 261.000 67.440 ;
      RECT 269.400 6.000 270.600 67.440 ;
    END
  END VDD
  OBS
    LAYER met1 ;
    RECT 0 0 281.060 73.440 ;
    LAYER met2 ;
    RECT 0 0 281.060 73.440 ;
    LAYER met3 ;
    RECT 0.800 0 281.060 73.440 ;
    RECT 0 0.000 0.800 5.850 ;
    RECT 0 6.150 0.800 6.450 ;
    RECT 0 6.750 0.800 7.050 ;
    RECT 0 7.350 0.800 7.650 ;
    RECT 0 7.950 0.800 8.250 ;
    RECT 0 8.550 0.800 8.850 ;
    RECT 0 9.150 0.800 9.450 ;
    RECT 0 9.750 0.800 10.050 ;
    RECT 0 10.350 0.800 10.650 ;
    RECT 0 10.950 0.800 11.250 ;
    RECT 0 11.550 0.800 11.850 ;
    RECT 0 12.150 0.800 12.450 ;
    RECT 0 12.750 0.800 13.050 ;
    RECT 0 13.350 0.800 13.650 ;
    RECT 0 13.950 0.800 14.250 ;
    RECT 0 14.550 0.800 21.450 ;
    RECT 0 21.750 0.800 22.050 ;
    RECT 0 22.350 0.800 22.650 ;
    RECT 0 22.950 0.800 23.250 ;
    RECT 0 23.550 0.800 23.850 ;
    RECT 0 24.150 0.800 24.450 ;
    RECT 0 24.750 0.800 25.050 ;
    RECT 0 25.350 0.800 25.650 ;
    RECT 0 25.950 0.800 26.250 ;
    RECT 0 26.550 0.800 26.850 ;
    RECT 0 27.150 0.800 27.450 ;
    RECT 0 27.750 0.800 28.050 ;
    RECT 0 28.350 0.800 28.650 ;
    RECT 0 28.950 0.800 29.250 ;
    RECT 0 29.550 0.800 29.850 ;
    RECT 0 30.150 0.800 37.050 ;
    RECT 0 37.350 0.800 37.650 ;
    RECT 0 37.950 0.800 38.250 ;
    RECT 0 38.550 0.800 38.850 ;
    RECT 0 39.150 0.800 39.450 ;
    RECT 0 39.750 0.800 40.050 ;
    RECT 0 40.350 0.800 40.650 ;
    RECT 0 40.950 0.800 41.250 ;
    RECT 0 41.550 0.800 41.850 ;
    RECT 0 42.150 0.800 42.450 ;
    RECT 0 42.750 0.800 43.050 ;
    RECT 0 43.350 0.800 43.650 ;
    RECT 0 43.950 0.800 44.250 ;
    RECT 0 44.550 0.800 44.850 ;
    RECT 0 45.150 0.800 45.450 ;
    RECT 0 45.750 0.800 52.650 ;
    RECT 0 52.950 0.800 53.250 ;
    RECT 0 53.550 0.800 53.850 ;
    RECT 0 54.150 0.800 54.450 ;
    RECT 0 54.750 0.800 55.050 ;
    RECT 0 55.350 0.800 55.650 ;
    RECT 0 55.950 0.800 62.850 ;
    RECT 0 63.150 0.800 63.450 ;
    RECT 0 63.750 0.800 64.050 ;
    RECT 0 64.350 0.800 73.440 ;
    LAYER met4 ;
    RECT 0 0 281.060 6.000 ;
    RECT 0 67.440 281.060 73.440 ;
    RECT 0.000 6.000 5.400 67.440 ;
    RECT 6.600 6.000 10.200 67.440 ;
    RECT 11.400 6.000 15.000 67.440 ;
    RECT 16.200 6.000 19.800 67.440 ;
    RECT 21.000 6.000 24.600 67.440 ;
    RECT 25.800 6.000 29.400 67.440 ;
    RECT 30.600 6.000 34.200 67.440 ;
    RECT 35.400 6.000 39.000 67.440 ;
    RECT 40.200 6.000 43.800 67.440 ;
    RECT 45.000 6.000 48.600 67.440 ;
    RECT 49.800 6.000 53.400 67.440 ;
    RECT 54.600 6.000 58.200 67.440 ;
    RECT 59.400 6.000 63.000 67.440 ;
    RECT 64.200 6.000 67.800 67.440 ;
    RECT 69.000 6.000 72.600 67.440 ;
    RECT 73.800 6.000 77.400 67.440 ;
    RECT 78.600 6.000 82.200 67.440 ;
    RECT 83.400 6.000 87.000 67.440 ;
    RECT 88.200 6.000 91.800 67.440 ;
    RECT 93.000 6.000 96.600 67.440 ;
    RECT 97.800 6.000 101.400 67.440 ;
    RECT 102.600 6.000 106.200 67.440 ;
    RECT 107.400 6.000 111.000 67.440 ;
    RECT 112.200 6.000 115.800 67.440 ;
    RECT 117.000 6.000 120.600 67.440 ;
    RECT 121.800 6.000 125.400 67.440 ;
    RECT 126.600 6.000 130.200 67.440 ;
    RECT 131.400 6.000 135.000 67.440 ;
    RECT 136.200 6.000 139.800 67.440 ;
    RECT 141.000 6.000 144.600 67.440 ;
    RECT 145.800 6.000 149.400 67.440 ;
    RECT 150.600 6.000 154.200 67.440 ;
    RECT 155.400 6.000 159.000 67.440 ;
    RECT 160.200 6.000 163.800 67.440 ;
    RECT 165.000 6.000 168.600 67.440 ;
    RECT 169.800 6.000 173.400 67.440 ;
    RECT 174.600 6.000 178.200 67.440 ;
    RECT 179.400 6.000 183.000 67.440 ;
    RECT 184.200 6.000 187.800 67.440 ;
    RECT 189.000 6.000 192.600 67.440 ;
    RECT 193.800 6.000 197.400 67.440 ;
    RECT 198.600 6.000 202.200 67.440 ;
    RECT 203.400 6.000 207.000 67.440 ;
    RECT 208.200 6.000 211.800 67.440 ;
    RECT 213.000 6.000 216.600 67.440 ;
    RECT 217.800 6.000 221.400 67.440 ;
    RECT 222.600 6.000 226.200 67.440 ;
    RECT 227.400 6.000 231.000 67.440 ;
    RECT 232.200 6.000 235.800 67.440 ;
    RECT 237.000 6.000 240.600 67.440 ;
    RECT 241.800 6.000 245.400 67.440 ;
    RECT 246.600 6.000 250.200 67.440 ;
    RECT 251.400 6.000 255.000 67.440 ;
    RECT 256.200 6.000 259.800 67.440 ;
    RECT 261.000 6.000 264.600 67.440 ;
    RECT 265.800 6.000 269.400 67.440 ;
    RECT 270.600 6.000 274.200 67.440 ;
    RECT 275.400 6.000 281.060 67.440 ;
    LAYER OVERLAP ;
    RECT 0 0 281.060 73.440 ;
  END
END fakeram130_64x15

END LIBRARY
