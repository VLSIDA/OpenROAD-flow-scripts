VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram130_2048x39
  FOREIGN fakeram130_2048x39 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 1031.320 BY 492.320 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 5.850 0.800 6.150 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 9.450 0.800 9.750 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 13.050 0.800 13.350 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 16.650 0.800 16.950 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 20.250 0.800 20.550 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 23.850 0.800 24.150 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 27.450 0.800 27.750 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 31.050 0.800 31.350 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 34.650 0.800 34.950 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 38.250 0.800 38.550 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 41.850 0.800 42.150 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 45.450 0.800 45.750 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 49.050 0.800 49.350 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 52.650 0.800 52.950 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 56.250 0.800 56.550 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 59.850 0.800 60.150 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 63.450 0.800 63.750 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 67.050 0.800 67.350 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 70.650 0.800 70.950 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 74.250 0.800 74.550 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 77.850 0.800 78.150 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 81.450 0.800 81.750 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 85.050 0.800 85.350 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 88.650 0.800 88.950 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 92.250 0.800 92.550 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 95.850 0.800 96.150 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 99.450 0.800 99.750 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 103.050 0.800 103.350 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 106.650 0.800 106.950 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 110.250 0.800 110.550 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 113.850 0.800 114.150 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 117.450 0.800 117.750 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 121.050 0.800 121.350 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 124.650 0.800 124.950 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 128.250 0.800 128.550 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 131.850 0.800 132.150 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 135.450 0.800 135.750 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 139.050 0.800 139.350 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 142.650 0.800 142.950 ;
    END
  END w_mask_in[38]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 144.450 0.800 144.750 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 148.050 0.800 148.350 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 151.650 0.800 151.950 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 155.250 0.800 155.550 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 158.850 0.800 159.150 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 162.450 0.800 162.750 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 166.050 0.800 166.350 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 169.650 0.800 169.950 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 173.250 0.800 173.550 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 176.850 0.800 177.150 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 180.450 0.800 180.750 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 184.050 0.800 184.350 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 187.650 0.800 187.950 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 191.250 0.800 191.550 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 194.850 0.800 195.150 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 198.450 0.800 198.750 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 202.050 0.800 202.350 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 205.650 0.800 205.950 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 209.250 0.800 209.550 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 212.850 0.800 213.150 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 216.450 0.800 216.750 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 220.050 0.800 220.350 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 223.650 0.800 223.950 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 227.250 0.800 227.550 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 230.850 0.800 231.150 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 234.450 0.800 234.750 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 238.050 0.800 238.350 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 241.650 0.800 241.950 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 245.250 0.800 245.550 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 248.850 0.800 249.150 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 252.450 0.800 252.750 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 256.050 0.800 256.350 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 259.650 0.800 259.950 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 263.250 0.800 263.550 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 266.850 0.800 267.150 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 270.450 0.800 270.750 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 274.050 0.800 274.350 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 277.650 0.800 277.950 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 281.250 0.800 281.550 ;
    END
  END rd_out[38]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 283.050 0.800 283.350 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 286.650 0.800 286.950 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 290.250 0.800 290.550 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 293.850 0.800 294.150 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 297.450 0.800 297.750 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 301.050 0.800 301.350 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 304.650 0.800 304.950 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 308.250 0.800 308.550 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 311.850 0.800 312.150 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 315.450 0.800 315.750 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 319.050 0.800 319.350 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 322.650 0.800 322.950 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 326.250 0.800 326.550 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 329.850 0.800 330.150 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 333.450 0.800 333.750 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 337.050 0.800 337.350 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 340.650 0.800 340.950 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 344.250 0.800 344.550 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 347.850 0.800 348.150 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 351.450 0.800 351.750 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 355.050 0.800 355.350 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 358.650 0.800 358.950 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 362.250 0.800 362.550 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 365.850 0.800 366.150 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 369.450 0.800 369.750 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 373.050 0.800 373.350 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 376.650 0.800 376.950 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 380.250 0.800 380.550 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 383.850 0.800 384.150 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 387.450 0.800 387.750 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 391.050 0.800 391.350 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 394.650 0.800 394.950 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 398.250 0.800 398.550 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 401.850 0.800 402.150 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 405.450 0.800 405.750 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 409.050 0.800 409.350 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 412.650 0.800 412.950 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 416.250 0.800 416.550 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 419.850 0.800 420.150 ;
    END
  END wd_in[38]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 421.650 0.800 421.950 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 425.250 0.800 425.550 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 428.850 0.800 429.150 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 432.450 0.800 432.750 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 436.050 0.800 436.350 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 439.650 0.800 439.950 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 443.250 0.800 443.550 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 446.850 0.800 447.150 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 450.450 0.800 450.750 ;
    END
  END addr_in[8]
  PIN addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 454.050 0.800 454.350 ;
    END
  END addr_in[9]
  PIN addr_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 457.650 0.800 457.950 ;
    END
  END addr_in[10]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 459.450 0.800 459.750 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 463.050 0.800 463.350 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 466.650 0.800 466.950 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
      RECT 5.400 6.000 6.600 486.320 ;
      RECT 15.000 6.000 16.200 486.320 ;
      RECT 24.600 6.000 25.800 486.320 ;
      RECT 34.200 6.000 35.400 486.320 ;
      RECT 43.800 6.000 45.000 486.320 ;
      RECT 53.400 6.000 54.600 486.320 ;
      RECT 63.000 6.000 64.200 486.320 ;
      RECT 72.600 6.000 73.800 486.320 ;
      RECT 82.200 6.000 83.400 486.320 ;
      RECT 91.800 6.000 93.000 486.320 ;
      RECT 101.400 6.000 102.600 486.320 ;
      RECT 111.000 6.000 112.200 486.320 ;
      RECT 120.600 6.000 121.800 486.320 ;
      RECT 130.200 6.000 131.400 486.320 ;
      RECT 139.800 6.000 141.000 486.320 ;
      RECT 149.400 6.000 150.600 486.320 ;
      RECT 159.000 6.000 160.200 486.320 ;
      RECT 168.600 6.000 169.800 486.320 ;
      RECT 178.200 6.000 179.400 486.320 ;
      RECT 187.800 6.000 189.000 486.320 ;
      RECT 197.400 6.000 198.600 486.320 ;
      RECT 207.000 6.000 208.200 486.320 ;
      RECT 216.600 6.000 217.800 486.320 ;
      RECT 226.200 6.000 227.400 486.320 ;
      RECT 235.800 6.000 237.000 486.320 ;
      RECT 245.400 6.000 246.600 486.320 ;
      RECT 255.000 6.000 256.200 486.320 ;
      RECT 264.600 6.000 265.800 486.320 ;
      RECT 274.200 6.000 275.400 486.320 ;
      RECT 283.800 6.000 285.000 486.320 ;
      RECT 293.400 6.000 294.600 486.320 ;
      RECT 303.000 6.000 304.200 486.320 ;
      RECT 312.600 6.000 313.800 486.320 ;
      RECT 322.200 6.000 323.400 486.320 ;
      RECT 331.800 6.000 333.000 486.320 ;
      RECT 341.400 6.000 342.600 486.320 ;
      RECT 351.000 6.000 352.200 486.320 ;
      RECT 360.600 6.000 361.800 486.320 ;
      RECT 370.200 6.000 371.400 486.320 ;
      RECT 379.800 6.000 381.000 486.320 ;
      RECT 389.400 6.000 390.600 486.320 ;
      RECT 399.000 6.000 400.200 486.320 ;
      RECT 408.600 6.000 409.800 486.320 ;
      RECT 418.200 6.000 419.400 486.320 ;
      RECT 427.800 6.000 429.000 486.320 ;
      RECT 437.400 6.000 438.600 486.320 ;
      RECT 447.000 6.000 448.200 486.320 ;
      RECT 456.600 6.000 457.800 486.320 ;
      RECT 466.200 6.000 467.400 486.320 ;
      RECT 475.800 6.000 477.000 486.320 ;
      RECT 485.400 6.000 486.600 486.320 ;
      RECT 495.000 6.000 496.200 486.320 ;
      RECT 504.600 6.000 505.800 486.320 ;
      RECT 514.200 6.000 515.400 486.320 ;
      RECT 523.800 6.000 525.000 486.320 ;
      RECT 533.400 6.000 534.600 486.320 ;
      RECT 543.000 6.000 544.200 486.320 ;
      RECT 552.600 6.000 553.800 486.320 ;
      RECT 562.200 6.000 563.400 486.320 ;
      RECT 571.800 6.000 573.000 486.320 ;
      RECT 581.400 6.000 582.600 486.320 ;
      RECT 591.000 6.000 592.200 486.320 ;
      RECT 600.600 6.000 601.800 486.320 ;
      RECT 610.200 6.000 611.400 486.320 ;
      RECT 619.800 6.000 621.000 486.320 ;
      RECT 629.400 6.000 630.600 486.320 ;
      RECT 639.000 6.000 640.200 486.320 ;
      RECT 648.600 6.000 649.800 486.320 ;
      RECT 658.200 6.000 659.400 486.320 ;
      RECT 667.800 6.000 669.000 486.320 ;
      RECT 677.400 6.000 678.600 486.320 ;
      RECT 687.000 6.000 688.200 486.320 ;
      RECT 696.600 6.000 697.800 486.320 ;
      RECT 706.200 6.000 707.400 486.320 ;
      RECT 715.800 6.000 717.000 486.320 ;
      RECT 725.400 6.000 726.600 486.320 ;
      RECT 735.000 6.000 736.200 486.320 ;
      RECT 744.600 6.000 745.800 486.320 ;
      RECT 754.200 6.000 755.400 486.320 ;
      RECT 763.800 6.000 765.000 486.320 ;
      RECT 773.400 6.000 774.600 486.320 ;
      RECT 783.000 6.000 784.200 486.320 ;
      RECT 792.600 6.000 793.800 486.320 ;
      RECT 802.200 6.000 803.400 486.320 ;
      RECT 811.800 6.000 813.000 486.320 ;
      RECT 821.400 6.000 822.600 486.320 ;
      RECT 831.000 6.000 832.200 486.320 ;
      RECT 840.600 6.000 841.800 486.320 ;
      RECT 850.200 6.000 851.400 486.320 ;
      RECT 859.800 6.000 861.000 486.320 ;
      RECT 869.400 6.000 870.600 486.320 ;
      RECT 879.000 6.000 880.200 486.320 ;
      RECT 888.600 6.000 889.800 486.320 ;
      RECT 898.200 6.000 899.400 486.320 ;
      RECT 907.800 6.000 909.000 486.320 ;
      RECT 917.400 6.000 918.600 486.320 ;
      RECT 927.000 6.000 928.200 486.320 ;
      RECT 936.600 6.000 937.800 486.320 ;
      RECT 946.200 6.000 947.400 486.320 ;
      RECT 955.800 6.000 957.000 486.320 ;
      RECT 965.400 6.000 966.600 486.320 ;
      RECT 975.000 6.000 976.200 486.320 ;
      RECT 984.600 6.000 985.800 486.320 ;
      RECT 994.200 6.000 995.400 486.320 ;
      RECT 1003.800 6.000 1005.000 486.320 ;
      RECT 1013.400 6.000 1014.600 486.320 ;
      RECT 1023.000 6.000 1024.200 486.320 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
      RECT 10.200 6.000 11.400 486.320 ;
      RECT 19.800 6.000 21.000 486.320 ;
      RECT 29.400 6.000 30.600 486.320 ;
      RECT 39.000 6.000 40.200 486.320 ;
      RECT 48.600 6.000 49.800 486.320 ;
      RECT 58.200 6.000 59.400 486.320 ;
      RECT 67.800 6.000 69.000 486.320 ;
      RECT 77.400 6.000 78.600 486.320 ;
      RECT 87.000 6.000 88.200 486.320 ;
      RECT 96.600 6.000 97.800 486.320 ;
      RECT 106.200 6.000 107.400 486.320 ;
      RECT 115.800 6.000 117.000 486.320 ;
      RECT 125.400 6.000 126.600 486.320 ;
      RECT 135.000 6.000 136.200 486.320 ;
      RECT 144.600 6.000 145.800 486.320 ;
      RECT 154.200 6.000 155.400 486.320 ;
      RECT 163.800 6.000 165.000 486.320 ;
      RECT 173.400 6.000 174.600 486.320 ;
      RECT 183.000 6.000 184.200 486.320 ;
      RECT 192.600 6.000 193.800 486.320 ;
      RECT 202.200 6.000 203.400 486.320 ;
      RECT 211.800 6.000 213.000 486.320 ;
      RECT 221.400 6.000 222.600 486.320 ;
      RECT 231.000 6.000 232.200 486.320 ;
      RECT 240.600 6.000 241.800 486.320 ;
      RECT 250.200 6.000 251.400 486.320 ;
      RECT 259.800 6.000 261.000 486.320 ;
      RECT 269.400 6.000 270.600 486.320 ;
      RECT 279.000 6.000 280.200 486.320 ;
      RECT 288.600 6.000 289.800 486.320 ;
      RECT 298.200 6.000 299.400 486.320 ;
      RECT 307.800 6.000 309.000 486.320 ;
      RECT 317.400 6.000 318.600 486.320 ;
      RECT 327.000 6.000 328.200 486.320 ;
      RECT 336.600 6.000 337.800 486.320 ;
      RECT 346.200 6.000 347.400 486.320 ;
      RECT 355.800 6.000 357.000 486.320 ;
      RECT 365.400 6.000 366.600 486.320 ;
      RECT 375.000 6.000 376.200 486.320 ;
      RECT 384.600 6.000 385.800 486.320 ;
      RECT 394.200 6.000 395.400 486.320 ;
      RECT 403.800 6.000 405.000 486.320 ;
      RECT 413.400 6.000 414.600 486.320 ;
      RECT 423.000 6.000 424.200 486.320 ;
      RECT 432.600 6.000 433.800 486.320 ;
      RECT 442.200 6.000 443.400 486.320 ;
      RECT 451.800 6.000 453.000 486.320 ;
      RECT 461.400 6.000 462.600 486.320 ;
      RECT 471.000 6.000 472.200 486.320 ;
      RECT 480.600 6.000 481.800 486.320 ;
      RECT 490.200 6.000 491.400 486.320 ;
      RECT 499.800 6.000 501.000 486.320 ;
      RECT 509.400 6.000 510.600 486.320 ;
      RECT 519.000 6.000 520.200 486.320 ;
      RECT 528.600 6.000 529.800 486.320 ;
      RECT 538.200 6.000 539.400 486.320 ;
      RECT 547.800 6.000 549.000 486.320 ;
      RECT 557.400 6.000 558.600 486.320 ;
      RECT 567.000 6.000 568.200 486.320 ;
      RECT 576.600 6.000 577.800 486.320 ;
      RECT 586.200 6.000 587.400 486.320 ;
      RECT 595.800 6.000 597.000 486.320 ;
      RECT 605.400 6.000 606.600 486.320 ;
      RECT 615.000 6.000 616.200 486.320 ;
      RECT 624.600 6.000 625.800 486.320 ;
      RECT 634.200 6.000 635.400 486.320 ;
      RECT 643.800 6.000 645.000 486.320 ;
      RECT 653.400 6.000 654.600 486.320 ;
      RECT 663.000 6.000 664.200 486.320 ;
      RECT 672.600 6.000 673.800 486.320 ;
      RECT 682.200 6.000 683.400 486.320 ;
      RECT 691.800 6.000 693.000 486.320 ;
      RECT 701.400 6.000 702.600 486.320 ;
      RECT 711.000 6.000 712.200 486.320 ;
      RECT 720.600 6.000 721.800 486.320 ;
      RECT 730.200 6.000 731.400 486.320 ;
      RECT 739.800 6.000 741.000 486.320 ;
      RECT 749.400 6.000 750.600 486.320 ;
      RECT 759.000 6.000 760.200 486.320 ;
      RECT 768.600 6.000 769.800 486.320 ;
      RECT 778.200 6.000 779.400 486.320 ;
      RECT 787.800 6.000 789.000 486.320 ;
      RECT 797.400 6.000 798.600 486.320 ;
      RECT 807.000 6.000 808.200 486.320 ;
      RECT 816.600 6.000 817.800 486.320 ;
      RECT 826.200 6.000 827.400 486.320 ;
      RECT 835.800 6.000 837.000 486.320 ;
      RECT 845.400 6.000 846.600 486.320 ;
      RECT 855.000 6.000 856.200 486.320 ;
      RECT 864.600 6.000 865.800 486.320 ;
      RECT 874.200 6.000 875.400 486.320 ;
      RECT 883.800 6.000 885.000 486.320 ;
      RECT 893.400 6.000 894.600 486.320 ;
      RECT 903.000 6.000 904.200 486.320 ;
      RECT 912.600 6.000 913.800 486.320 ;
      RECT 922.200 6.000 923.400 486.320 ;
      RECT 931.800 6.000 933.000 486.320 ;
      RECT 941.400 6.000 942.600 486.320 ;
      RECT 951.000 6.000 952.200 486.320 ;
      RECT 960.600 6.000 961.800 486.320 ;
      RECT 970.200 6.000 971.400 486.320 ;
      RECT 979.800 6.000 981.000 486.320 ;
      RECT 989.400 6.000 990.600 486.320 ;
      RECT 999.000 6.000 1000.200 486.320 ;
      RECT 1008.600 6.000 1009.800 486.320 ;
      RECT 1018.200 6.000 1019.400 486.320 ;
    END
  END VDD
  OBS
    LAYER met1 ;
    RECT 0 0 1031.320 492.320 ;
    LAYER met2 ;
    RECT 0 0 1031.320 492.320 ;
    LAYER met3 ;
    RECT 0.800 0 1031.320 492.320 ;
    RECT 0 0.000 0.800 5.850 ;
    RECT 0 6.150 0.800 9.450 ;
    RECT 0 9.750 0.800 13.050 ;
    RECT 0 13.350 0.800 16.650 ;
    RECT 0 16.950 0.800 20.250 ;
    RECT 0 20.550 0.800 23.850 ;
    RECT 0 24.150 0.800 27.450 ;
    RECT 0 27.750 0.800 31.050 ;
    RECT 0 31.350 0.800 34.650 ;
    RECT 0 34.950 0.800 38.250 ;
    RECT 0 38.550 0.800 41.850 ;
    RECT 0 42.150 0.800 45.450 ;
    RECT 0 45.750 0.800 49.050 ;
    RECT 0 49.350 0.800 52.650 ;
    RECT 0 52.950 0.800 56.250 ;
    RECT 0 56.550 0.800 59.850 ;
    RECT 0 60.150 0.800 63.450 ;
    RECT 0 63.750 0.800 67.050 ;
    RECT 0 67.350 0.800 70.650 ;
    RECT 0 70.950 0.800 74.250 ;
    RECT 0 74.550 0.800 77.850 ;
    RECT 0 78.150 0.800 81.450 ;
    RECT 0 81.750 0.800 85.050 ;
    RECT 0 85.350 0.800 88.650 ;
    RECT 0 88.950 0.800 92.250 ;
    RECT 0 92.550 0.800 95.850 ;
    RECT 0 96.150 0.800 99.450 ;
    RECT 0 99.750 0.800 103.050 ;
    RECT 0 103.350 0.800 106.650 ;
    RECT 0 106.950 0.800 110.250 ;
    RECT 0 110.550 0.800 113.850 ;
    RECT 0 114.150 0.800 117.450 ;
    RECT 0 117.750 0.800 121.050 ;
    RECT 0 121.350 0.800 124.650 ;
    RECT 0 124.950 0.800 128.250 ;
    RECT 0 128.550 0.800 131.850 ;
    RECT 0 132.150 0.800 135.450 ;
    RECT 0 135.750 0.800 139.050 ;
    RECT 0 139.350 0.800 142.650 ;
    RECT 0 142.950 0.800 144.450 ;
    RECT 0 144.750 0.800 148.050 ;
    RECT 0 148.350 0.800 151.650 ;
    RECT 0 151.950 0.800 155.250 ;
    RECT 0 155.550 0.800 158.850 ;
    RECT 0 159.150 0.800 162.450 ;
    RECT 0 162.750 0.800 166.050 ;
    RECT 0 166.350 0.800 169.650 ;
    RECT 0 169.950 0.800 173.250 ;
    RECT 0 173.550 0.800 176.850 ;
    RECT 0 177.150 0.800 180.450 ;
    RECT 0 180.750 0.800 184.050 ;
    RECT 0 184.350 0.800 187.650 ;
    RECT 0 187.950 0.800 191.250 ;
    RECT 0 191.550 0.800 194.850 ;
    RECT 0 195.150 0.800 198.450 ;
    RECT 0 198.750 0.800 202.050 ;
    RECT 0 202.350 0.800 205.650 ;
    RECT 0 205.950 0.800 209.250 ;
    RECT 0 209.550 0.800 212.850 ;
    RECT 0 213.150 0.800 216.450 ;
    RECT 0 216.750 0.800 220.050 ;
    RECT 0 220.350 0.800 223.650 ;
    RECT 0 223.950 0.800 227.250 ;
    RECT 0 227.550 0.800 230.850 ;
    RECT 0 231.150 0.800 234.450 ;
    RECT 0 234.750 0.800 238.050 ;
    RECT 0 238.350 0.800 241.650 ;
    RECT 0 241.950 0.800 245.250 ;
    RECT 0 245.550 0.800 248.850 ;
    RECT 0 249.150 0.800 252.450 ;
    RECT 0 252.750 0.800 256.050 ;
    RECT 0 256.350 0.800 259.650 ;
    RECT 0 259.950 0.800 263.250 ;
    RECT 0 263.550 0.800 266.850 ;
    RECT 0 267.150 0.800 270.450 ;
    RECT 0 270.750 0.800 274.050 ;
    RECT 0 274.350 0.800 277.650 ;
    RECT 0 277.950 0.800 281.250 ;
    RECT 0 281.550 0.800 283.050 ;
    RECT 0 283.350 0.800 286.650 ;
    RECT 0 286.950 0.800 290.250 ;
    RECT 0 290.550 0.800 293.850 ;
    RECT 0 294.150 0.800 297.450 ;
    RECT 0 297.750 0.800 301.050 ;
    RECT 0 301.350 0.800 304.650 ;
    RECT 0 304.950 0.800 308.250 ;
    RECT 0 308.550 0.800 311.850 ;
    RECT 0 312.150 0.800 315.450 ;
    RECT 0 315.750 0.800 319.050 ;
    RECT 0 319.350 0.800 322.650 ;
    RECT 0 322.950 0.800 326.250 ;
    RECT 0 326.550 0.800 329.850 ;
    RECT 0 330.150 0.800 333.450 ;
    RECT 0 333.750 0.800 337.050 ;
    RECT 0 337.350 0.800 340.650 ;
    RECT 0 340.950 0.800 344.250 ;
    RECT 0 344.550 0.800 347.850 ;
    RECT 0 348.150 0.800 351.450 ;
    RECT 0 351.750 0.800 355.050 ;
    RECT 0 355.350 0.800 358.650 ;
    RECT 0 358.950 0.800 362.250 ;
    RECT 0 362.550 0.800 365.850 ;
    RECT 0 366.150 0.800 369.450 ;
    RECT 0 369.750 0.800 373.050 ;
    RECT 0 373.350 0.800 376.650 ;
    RECT 0 376.950 0.800 380.250 ;
    RECT 0 380.550 0.800 383.850 ;
    RECT 0 384.150 0.800 387.450 ;
    RECT 0 387.750 0.800 391.050 ;
    RECT 0 391.350 0.800 394.650 ;
    RECT 0 394.950 0.800 398.250 ;
    RECT 0 398.550 0.800 401.850 ;
    RECT 0 402.150 0.800 405.450 ;
    RECT 0 405.750 0.800 409.050 ;
    RECT 0 409.350 0.800 412.650 ;
    RECT 0 412.950 0.800 416.250 ;
    RECT 0 416.550 0.800 419.850 ;
    RECT 0 420.150 0.800 421.650 ;
    RECT 0 421.950 0.800 425.250 ;
    RECT 0 425.550 0.800 428.850 ;
    RECT 0 429.150 0.800 432.450 ;
    RECT 0 432.750 0.800 436.050 ;
    RECT 0 436.350 0.800 439.650 ;
    RECT 0 439.950 0.800 443.250 ;
    RECT 0 443.550 0.800 446.850 ;
    RECT 0 447.150 0.800 450.450 ;
    RECT 0 450.750 0.800 454.050 ;
    RECT 0 454.350 0.800 457.650 ;
    RECT 0 457.950 0.800 459.450 ;
    RECT 0 459.750 0.800 463.050 ;
    RECT 0 463.350 0.800 466.650 ;
    RECT 0 466.950 0.800 492.320 ;
    LAYER met4 ;
    RECT 0 0 1031.320 6.000 ;
    RECT 0 486.320 1031.320 492.320 ;
    RECT 0.000 6.000 5.400 486.320 ;
    RECT 6.600 6.000 10.200 486.320 ;
    RECT 11.400 6.000 15.000 486.320 ;
    RECT 16.200 6.000 19.800 486.320 ;
    RECT 21.000 6.000 24.600 486.320 ;
    RECT 25.800 6.000 29.400 486.320 ;
    RECT 30.600 6.000 34.200 486.320 ;
    RECT 35.400 6.000 39.000 486.320 ;
    RECT 40.200 6.000 43.800 486.320 ;
    RECT 45.000 6.000 48.600 486.320 ;
    RECT 49.800 6.000 53.400 486.320 ;
    RECT 54.600 6.000 58.200 486.320 ;
    RECT 59.400 6.000 63.000 486.320 ;
    RECT 64.200 6.000 67.800 486.320 ;
    RECT 69.000 6.000 72.600 486.320 ;
    RECT 73.800 6.000 77.400 486.320 ;
    RECT 78.600 6.000 82.200 486.320 ;
    RECT 83.400 6.000 87.000 486.320 ;
    RECT 88.200 6.000 91.800 486.320 ;
    RECT 93.000 6.000 96.600 486.320 ;
    RECT 97.800 6.000 101.400 486.320 ;
    RECT 102.600 6.000 106.200 486.320 ;
    RECT 107.400 6.000 111.000 486.320 ;
    RECT 112.200 6.000 115.800 486.320 ;
    RECT 117.000 6.000 120.600 486.320 ;
    RECT 121.800 6.000 125.400 486.320 ;
    RECT 126.600 6.000 130.200 486.320 ;
    RECT 131.400 6.000 135.000 486.320 ;
    RECT 136.200 6.000 139.800 486.320 ;
    RECT 141.000 6.000 144.600 486.320 ;
    RECT 145.800 6.000 149.400 486.320 ;
    RECT 150.600 6.000 154.200 486.320 ;
    RECT 155.400 6.000 159.000 486.320 ;
    RECT 160.200 6.000 163.800 486.320 ;
    RECT 165.000 6.000 168.600 486.320 ;
    RECT 169.800 6.000 173.400 486.320 ;
    RECT 174.600 6.000 178.200 486.320 ;
    RECT 179.400 6.000 183.000 486.320 ;
    RECT 184.200 6.000 187.800 486.320 ;
    RECT 189.000 6.000 192.600 486.320 ;
    RECT 193.800 6.000 197.400 486.320 ;
    RECT 198.600 6.000 202.200 486.320 ;
    RECT 203.400 6.000 207.000 486.320 ;
    RECT 208.200 6.000 211.800 486.320 ;
    RECT 213.000 6.000 216.600 486.320 ;
    RECT 217.800 6.000 221.400 486.320 ;
    RECT 222.600 6.000 226.200 486.320 ;
    RECT 227.400 6.000 231.000 486.320 ;
    RECT 232.200 6.000 235.800 486.320 ;
    RECT 237.000 6.000 240.600 486.320 ;
    RECT 241.800 6.000 245.400 486.320 ;
    RECT 246.600 6.000 250.200 486.320 ;
    RECT 251.400 6.000 255.000 486.320 ;
    RECT 256.200 6.000 259.800 486.320 ;
    RECT 261.000 6.000 264.600 486.320 ;
    RECT 265.800 6.000 269.400 486.320 ;
    RECT 270.600 6.000 274.200 486.320 ;
    RECT 275.400 6.000 279.000 486.320 ;
    RECT 280.200 6.000 283.800 486.320 ;
    RECT 285.000 6.000 288.600 486.320 ;
    RECT 289.800 6.000 293.400 486.320 ;
    RECT 294.600 6.000 298.200 486.320 ;
    RECT 299.400 6.000 303.000 486.320 ;
    RECT 304.200 6.000 307.800 486.320 ;
    RECT 309.000 6.000 312.600 486.320 ;
    RECT 313.800 6.000 317.400 486.320 ;
    RECT 318.600 6.000 322.200 486.320 ;
    RECT 323.400 6.000 327.000 486.320 ;
    RECT 328.200 6.000 331.800 486.320 ;
    RECT 333.000 6.000 336.600 486.320 ;
    RECT 337.800 6.000 341.400 486.320 ;
    RECT 342.600 6.000 346.200 486.320 ;
    RECT 347.400 6.000 351.000 486.320 ;
    RECT 352.200 6.000 355.800 486.320 ;
    RECT 357.000 6.000 360.600 486.320 ;
    RECT 361.800 6.000 365.400 486.320 ;
    RECT 366.600 6.000 370.200 486.320 ;
    RECT 371.400 6.000 375.000 486.320 ;
    RECT 376.200 6.000 379.800 486.320 ;
    RECT 381.000 6.000 384.600 486.320 ;
    RECT 385.800 6.000 389.400 486.320 ;
    RECT 390.600 6.000 394.200 486.320 ;
    RECT 395.400 6.000 399.000 486.320 ;
    RECT 400.200 6.000 403.800 486.320 ;
    RECT 405.000 6.000 408.600 486.320 ;
    RECT 409.800 6.000 413.400 486.320 ;
    RECT 414.600 6.000 418.200 486.320 ;
    RECT 419.400 6.000 423.000 486.320 ;
    RECT 424.200 6.000 427.800 486.320 ;
    RECT 429.000 6.000 432.600 486.320 ;
    RECT 433.800 6.000 437.400 486.320 ;
    RECT 438.600 6.000 442.200 486.320 ;
    RECT 443.400 6.000 447.000 486.320 ;
    RECT 448.200 6.000 451.800 486.320 ;
    RECT 453.000 6.000 456.600 486.320 ;
    RECT 457.800 6.000 461.400 486.320 ;
    RECT 462.600 6.000 466.200 486.320 ;
    RECT 467.400 6.000 471.000 486.320 ;
    RECT 472.200 6.000 475.800 486.320 ;
    RECT 477.000 6.000 480.600 486.320 ;
    RECT 481.800 6.000 485.400 486.320 ;
    RECT 486.600 6.000 490.200 486.320 ;
    RECT 491.400 6.000 495.000 486.320 ;
    RECT 496.200 6.000 499.800 486.320 ;
    RECT 501.000 6.000 504.600 486.320 ;
    RECT 505.800 6.000 509.400 486.320 ;
    RECT 510.600 6.000 514.200 486.320 ;
    RECT 515.400 6.000 519.000 486.320 ;
    RECT 520.200 6.000 523.800 486.320 ;
    RECT 525.000 6.000 528.600 486.320 ;
    RECT 529.800 6.000 533.400 486.320 ;
    RECT 534.600 6.000 538.200 486.320 ;
    RECT 539.400 6.000 543.000 486.320 ;
    RECT 544.200 6.000 547.800 486.320 ;
    RECT 549.000 6.000 552.600 486.320 ;
    RECT 553.800 6.000 557.400 486.320 ;
    RECT 558.600 6.000 562.200 486.320 ;
    RECT 563.400 6.000 567.000 486.320 ;
    RECT 568.200 6.000 571.800 486.320 ;
    RECT 573.000 6.000 576.600 486.320 ;
    RECT 577.800 6.000 581.400 486.320 ;
    RECT 582.600 6.000 586.200 486.320 ;
    RECT 587.400 6.000 591.000 486.320 ;
    RECT 592.200 6.000 595.800 486.320 ;
    RECT 597.000 6.000 600.600 486.320 ;
    RECT 601.800 6.000 605.400 486.320 ;
    RECT 606.600 6.000 610.200 486.320 ;
    RECT 611.400 6.000 615.000 486.320 ;
    RECT 616.200 6.000 619.800 486.320 ;
    RECT 621.000 6.000 624.600 486.320 ;
    RECT 625.800 6.000 629.400 486.320 ;
    RECT 630.600 6.000 634.200 486.320 ;
    RECT 635.400 6.000 639.000 486.320 ;
    RECT 640.200 6.000 643.800 486.320 ;
    RECT 645.000 6.000 648.600 486.320 ;
    RECT 649.800 6.000 653.400 486.320 ;
    RECT 654.600 6.000 658.200 486.320 ;
    RECT 659.400 6.000 663.000 486.320 ;
    RECT 664.200 6.000 667.800 486.320 ;
    RECT 669.000 6.000 672.600 486.320 ;
    RECT 673.800 6.000 677.400 486.320 ;
    RECT 678.600 6.000 682.200 486.320 ;
    RECT 683.400 6.000 687.000 486.320 ;
    RECT 688.200 6.000 691.800 486.320 ;
    RECT 693.000 6.000 696.600 486.320 ;
    RECT 697.800 6.000 701.400 486.320 ;
    RECT 702.600 6.000 706.200 486.320 ;
    RECT 707.400 6.000 711.000 486.320 ;
    RECT 712.200 6.000 715.800 486.320 ;
    RECT 717.000 6.000 720.600 486.320 ;
    RECT 721.800 6.000 725.400 486.320 ;
    RECT 726.600 6.000 730.200 486.320 ;
    RECT 731.400 6.000 735.000 486.320 ;
    RECT 736.200 6.000 739.800 486.320 ;
    RECT 741.000 6.000 744.600 486.320 ;
    RECT 745.800 6.000 749.400 486.320 ;
    RECT 750.600 6.000 754.200 486.320 ;
    RECT 755.400 6.000 759.000 486.320 ;
    RECT 760.200 6.000 763.800 486.320 ;
    RECT 765.000 6.000 768.600 486.320 ;
    RECT 769.800 6.000 773.400 486.320 ;
    RECT 774.600 6.000 778.200 486.320 ;
    RECT 779.400 6.000 783.000 486.320 ;
    RECT 784.200 6.000 787.800 486.320 ;
    RECT 789.000 6.000 792.600 486.320 ;
    RECT 793.800 6.000 797.400 486.320 ;
    RECT 798.600 6.000 802.200 486.320 ;
    RECT 803.400 6.000 807.000 486.320 ;
    RECT 808.200 6.000 811.800 486.320 ;
    RECT 813.000 6.000 816.600 486.320 ;
    RECT 817.800 6.000 821.400 486.320 ;
    RECT 822.600 6.000 826.200 486.320 ;
    RECT 827.400 6.000 831.000 486.320 ;
    RECT 832.200 6.000 835.800 486.320 ;
    RECT 837.000 6.000 840.600 486.320 ;
    RECT 841.800 6.000 845.400 486.320 ;
    RECT 846.600 6.000 850.200 486.320 ;
    RECT 851.400 6.000 855.000 486.320 ;
    RECT 856.200 6.000 859.800 486.320 ;
    RECT 861.000 6.000 864.600 486.320 ;
    RECT 865.800 6.000 869.400 486.320 ;
    RECT 870.600 6.000 874.200 486.320 ;
    RECT 875.400 6.000 879.000 486.320 ;
    RECT 880.200 6.000 883.800 486.320 ;
    RECT 885.000 6.000 888.600 486.320 ;
    RECT 889.800 6.000 893.400 486.320 ;
    RECT 894.600 6.000 898.200 486.320 ;
    RECT 899.400 6.000 903.000 486.320 ;
    RECT 904.200 6.000 907.800 486.320 ;
    RECT 909.000 6.000 912.600 486.320 ;
    RECT 913.800 6.000 917.400 486.320 ;
    RECT 918.600 6.000 922.200 486.320 ;
    RECT 923.400 6.000 927.000 486.320 ;
    RECT 928.200 6.000 931.800 486.320 ;
    RECT 933.000 6.000 936.600 486.320 ;
    RECT 937.800 6.000 941.400 486.320 ;
    RECT 942.600 6.000 946.200 486.320 ;
    RECT 947.400 6.000 951.000 486.320 ;
    RECT 952.200 6.000 955.800 486.320 ;
    RECT 957.000 6.000 960.600 486.320 ;
    RECT 961.800 6.000 965.400 486.320 ;
    RECT 966.600 6.000 970.200 486.320 ;
    RECT 971.400 6.000 975.000 486.320 ;
    RECT 976.200 6.000 979.800 486.320 ;
    RECT 981.000 6.000 984.600 486.320 ;
    RECT 985.800 6.000 989.400 486.320 ;
    RECT 990.600 6.000 994.200 486.320 ;
    RECT 995.400 6.000 999.000 486.320 ;
    RECT 1000.200 6.000 1003.800 486.320 ;
    RECT 1005.000 6.000 1008.600 486.320 ;
    RECT 1009.800 6.000 1013.400 486.320 ;
    RECT 1014.600 6.000 1018.200 486.320 ;
    RECT 1019.400 6.000 1023.000 486.320 ;
    RECT 1024.200 6.000 1031.320 486.320 ;
    LAYER OVERLAP ;
    RECT 0 0 1031.320 492.320 ;
  END
END fakeram130_2048x39

END LIBRARY
